�        �B��  �1��м |PP��|f`fh    fh   f�|f�|f�   f�   f��f1�f�   f��RVf�6|f�6|PRh h �|����^Zf�>|�uf�|f�|f��   �faf�                                                                                                                                                                                                                                                                                                                                                                         U��,��������������        ��   �� ��   ��    ��  �м PP�� ���f`fh    fh	   f�|f�|f� 0 f��   f��f1�f�   f��RVf�6|f�6|PRh h �|���sm^Zf�>|�uf�|f�|f��   �fafPfSfWj �f1�&f� &f�E   f� �  f�   f�PAMS���f�� u�f_f[fX(��p��p �"�f�   f� �؎���f���м   �    �   �   ��    �   �   �  �   ����   �  �   �   �   ���   "� �   �"�� 0 �  ���  � ����V��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �!  ���U��PQRSTUVW1ҋE�    f����E��} u����Ӊ_^]\[ZYX�� U��QRSTUVW1ҋE�    f����E���rh    X_^]\[ZY�� h   X_^]\[ZY�� U��R�E�U��rh    XZ�� h   XZ�� �U��PQRSTUVW�u�}�M�_^]\[ZYX�� U��PQRSTUVW�u�}�M�f�_^]\[ZYX�� ���U��PQRSTUVW�}�U�������������ЋU�����у��_^]\[ZYX�� �U��PQRSTUVW�}�Uf����f�ЋU�����у��f�_^]\[ZYX�� �U��PQRSTUVW�}�E�M�_^]\[ZYX�� ��0<9~�U��PQRSTUVW�]�u�   ������������F��$������F����� _^]\[ZYX�� U��PQRSTUVW�E�u1ɻ
   1����0RA��u�Z�F��� _^]\[ZYX��  �   U��P�E��E��� h�  P�5�������X�� U��PQRSTUVW�E�P   f��Ef�!�������f���f�_^]\[ZYX�� U��PQRSTUVW1ɋM��M��M�E�P   f��E����f�_^]\[ZYX�� PQRSTUVW�5�����Ơ   �   jPVW��������Ơ   ��=����   �G�0�jPPW�*���_^]\[ZYX�                                                
 U���u�u������u�@���u�D���8��    �<��    �5<���58�������� �<���8��    �=<��v�����<��   �5<���58������Ã=8�� vC�8���5@���5D���  h����$   �D���@���8���5<���58���2����U��PQRSTUVW�u1��< u_^]\[ZYX�� <
u�O����@<u�~����5�5<���58���5D���5@��P�����8���5<���58��������_^]\[ZYX��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ����U��PQRSTUVW���E������]�Mf���f�Xf�@ �@ �H�_^]\[ZYX�� P�p$�p�X�P� � XP� �X�RESET SYSTEM! jj�H����5@���5D���Yexc - 0,  Fault. #DE - Divide Error Exception. Induced (div, idiv). Induced (div, idiv). h������hH�������D���@���5@���5D��h����{����D���@�����jj�����5@���5D���-exc - 1,  Fault/Trap. #DB - Debug Exception. h�������hH�������D���@���5@���5D��h���������D���@�����jj�
����5@���5D���Cexc - 2,  Interrupt. Hardware failure. Induced (Hardware failure). hN������hH���u����D���@���5@���5D��h����S����D���@�����jj�k����5@���5D���=exc - 3,  Trap. #BP - Breakpoint Exception. Induced (int 3). h��������hH��������D���@���jj������5@���5D���:exc - 4,  Trap. #OF - Overflow Exception. Induced (into). hb���t���hH���j����D���@���jj�����5@���5D���Hexc - 5,  Fault. #BR - BOUND Range Exceeded Exception. Induced (bound). h��������hH��������D���@���5@���5D��h���������D���@�����jj������5@���5D���Lexc - 6,  Fault. #UD - Invalid Opcode Exception. Induced (invalid command). hx���L���hH���B����D���@���5@���5D��h���� ����D���@�����jj�8����5@���5D���Lexc - 7,  Fault. #NM - Device Not Available Exception. Induced (esc, wait). h ������hH�������D���@���5@���5D��h����x����D���@�����jj�����5@���5D���/exc - 8,  Abort. #DF - Double Fault Exception. h�������hH�������D���@���5@���5D��h���������D���@�����jj�����5@���5D���8exc - 9,  Fault. The output of the coprocessor segment. hS������hH���{����D���@���5@���5D��h����Y����D���@�����Xjj�p����5@���5D���Texc - 10, Fault. #TS - Invalid TSS Exception. Induced (jmp, call, iret, interrupt). h���������D���@���5@���5D���Error:  h`�������D���@���5@���5D���@��   h��P�D���h���q����D���@���5@���5D��h����O����D���@�����Xjj�f����5@���5D���Uexc - 11, Fault. #NP - Segment Not Present. Induced (segment register load command). h��������hH�������D���@���5@���5D���Error:  hu�������D���@���5@���5D���@��   h��P�/���h���\����D���@���5@���5D��h����:����D���@�����Xjj�Q����5@���5D���nexc - 12, Fault. #SS - Stack Fault Exception. Induced (stack access command). Induced (stack access command). h������hH�������D���@���5@���5D���Error:  h����e����D���@���5@���5D���@��   h��P����h���.����D���@���5@���5D��h��������D���@�����Xjj�#����5@���5D���Vexc - 13, Fault. #GP - General Protection Exception. Induced (memory access command). h5������hH���{����D���@���5@���5D���Error:  h����O����D���@���5@���5D���@��   h��P�����h�������D���@���5@���5D��h���������D���@�����[jj�����5@���5D���-exc - 14, Fault. #PF - Page-Fault Exception. hK������hH�������D���@���5@���5D���0Induced (memory access command). Page addres =  h����:����D���@�� ��5@���5D���@��   h��P����h��� ����D���@���5@���5D���@��   �h h>�������hH��������D���@���5@���5D���Error code -  hn�������D���@���5@���5D���@��   h��S�����h���]����D���@���5@���5D���@��   �h h����-���hH���#����D���@��j S������u=�5@���5D���Page present h�������hH��������D���@���?�5@���5D���Page not present h[������hH�������D���@��jS�������u;�5@���5D���Write page h����^���hH���T����D���@���8�5@���5D���
Read page h����$���hH�������D���@��jS�v�����u:�5@���5D���
User mode h'�������hH��������D���@���:�5@���5D���Kernel mode ha������hH�������D���@��jS�������uD�5@���5D���Write reserved bits h����T���hH���J����D���@���0�5@���5D���- h����"���hH�������D���@��jS�t�����uA�5@���5D���Read instruction h)�������hH��������D���@���0�5@���5D���- hj������hH�������D���@���5@���5D��h����x����D���@�����jj�����5@���5D���Shit!!! h����@���hH���6����D���@���5@���5D��h��������D���@�����jj�,����5@���5D���Jexc - 16, Fault. #MF - x87 FPU Floating-Point Error. Induced (esc, wait). h,������hH�������D���@���5@���5D��h����n����D���@�����Xjj�����5@���5D���sexc - 17, Fault. #AC - Alignment Check Exception.Induced (memory access command). Induced (memory access command). h���������D���@���5@���5D���Error:  hj�������D���@���5@���5D���@��   h��P�:���h���g����D���@���5@���5D��h����E����D���@�����            QRSTUVW1ҹ    Rh  ���;����� u
RX_^]\[ZY�B��h    X_^]\[ZYÐ��PQRSTUVW�=���   sKjj�����5@���5D���Not free memory! hW������hH�������D���@������`���jPh  ���k������-���   _^]\[ZYXÐU��PQRSTUVW�M�E��j Ph  ���3�������   �E   ��_^]\[ZYX��    �    ����        ��   �� ��   ��   ����PQRSTUVW��`h   j�h  ���/�������  ����   �������������Q�5����@���a �% �������_^]\[ZYXÐU��PQRSTUVW� �����
���E����   = ���_^]\[ZYX�� ��U��PQRSTUVW�M�u���}��
��������� u�:������������% ���P�����EE�� ���}�E   �_^]\[ZYX�� �    `��0 ���P� � XP� �Xa�                        �`�1��`�=_ ��r
�_ ��    �=_ ����K ���_ ���aP�a4P�a�P� � XP� �Xa���5@���5D��V�_����D���@���ϐ��  1234567890-= qwertyuiop[]
 asdfghjkl;'` \zxcvbnm,./ *                  -   +                              ���  !@#$%^&*()_+ QWERTYUIOP{}
 ASDFGHJKL:"~ |ZXCVBNM<>? *                  -   +                               Ph � ���f�c  f�!��Xj�@��j �D���5D���5@���f����    P�� XP� �!XP��!XP��!XP���!XP��XP�(�XP��XP��XP���Xh�  j h��������h�   h���j �K���h�   h���j!�:���j j j"�/���h�   h���j#����h�   h���j$����h�   h���j%�����h�   h���j&�����h�   h���j'�����h�   h���j(�����h�   h���j)����h�   h���j*����h�   h���j+����h�   h���j,����h�   h���j-�t���h�   h���j.�c���h�   h���j/�R������h�   h���j �:���h�   h���j�)���h�   h7��j����h�   h���j����h�   hK��j�����h�   h���j�����h�   ha��j�����h�   h	��j�����h�   h���j����h�   h<��j	����h�   h���j
����h�   h���j����h�   h���j�n���h�   h��j�]���h�   h3��j�L���h�   h���j�;���h�   h��j�*���h�   h���j��������Ph�   h4 ��j ����P�6�CX��.  P���@XP���@XXh�   hd ��j!�����h�   h� ��j0����������5@���5D���@��   �$Velcome to Varania OS! version: 1.0 h�$������hH��������D���@�������jjPh   ����jhX%��h   �`�����?����`%���0�Prg1
Hello
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             